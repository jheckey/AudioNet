/* 8-bit Grey-code decoder
Copyright: Hectic Tech, 2012, all rights reserved
Author: Jeff Heckey (jheckey@gmail.com)

Module: gc2bin8

Purpose: 
    Decodes Grey-coded to binary

Function:
    Decodes Grey-coded bytes to binary
*/

module gc2bin8 (
    input  wire [7:0]  gc,
    output wire [7:0]  bin
);

reg  [7:0]     bin_r;

assign bin = bin_r;

always @* begin
    case (gc)
        8'b00000000: bin_r = 8'b00000000;  // gc: 0, bin: 0
        8'b00000001: bin_r = 8'b00000001;  // gc: 1, bin: 1
        8'b00000011: bin_r = 8'b00000010;  // gc: 3, bin: 2
        8'b00000010: bin_r = 8'b00000011;  // gc: 2, bin: 3
        8'b00000110: bin_r = 8'b00000100;  // gc: 6, bin: 4
        8'b00000111: bin_r = 8'b00000101;  // gc: 7, bin: 5
        8'b00000101: bin_r = 8'b00000110;  // gc: 5, bin: 6
        8'b00000100: bin_r = 8'b00000111;  // gc: 4, bin: 7
        8'b00001100: bin_r = 8'b00001000;  // gc: 12, bin: 8
        8'b00001101: bin_r = 8'b00001001;  // gc: 13, bin: 9
        8'b00001111: bin_r = 8'b00001010;  // gc: 15, bin: 10
        8'b00001110: bin_r = 8'b00001011;  // gc: 14, bin: 11
        8'b00001010: bin_r = 8'b00001100;  // gc: 10, bin: 12
        8'b00001011: bin_r = 8'b00001101;  // gc: 11, bin: 13
        8'b00001001: bin_r = 8'b00001110;  // gc: 9, bin: 14
        8'b00001000: bin_r = 8'b00001111;  // gc: 8, bin: 15
        8'b00011000: bin_r = 8'b00010000;  // gc: 24, bin: 16
        8'b00011001: bin_r = 8'b00010001;  // gc: 25, bin: 17
        8'b00011011: bin_r = 8'b00010010;  // gc: 27, bin: 18
        8'b00011010: bin_r = 8'b00010011;  // gc: 26, bin: 19
        8'b00011110: bin_r = 8'b00010100;  // gc: 30, bin: 20
        8'b00011111: bin_r = 8'b00010101;  // gc: 31, bin: 21
        8'b00011101: bin_r = 8'b00010110;  // gc: 29, bin: 22
        8'b00011100: bin_r = 8'b00010111;  // gc: 28, bin: 23
        8'b00010100: bin_r = 8'b00011000;  // gc: 20, bin: 24
        8'b00010101: bin_r = 8'b00011001;  // gc: 21, bin: 25
        8'b00010111: bin_r = 8'b00011010;  // gc: 23, bin: 26
        8'b00010110: bin_r = 8'b00011011;  // gc: 22, bin: 27
        8'b00010010: bin_r = 8'b00011100;  // gc: 18, bin: 28
        8'b00010011: bin_r = 8'b00011101;  // gc: 19, bin: 29
        8'b00010001: bin_r = 8'b00011110;  // gc: 17, bin: 30
        8'b00010000: bin_r = 8'b00011111;  // gc: 16, bin: 31
        8'b00110000: bin_r = 8'b00100000;  // gc: 48, bin: 32
        8'b00110001: bin_r = 8'b00100001;  // gc: 49, bin: 33
        8'b00110011: bin_r = 8'b00100010;  // gc: 51, bin: 34
        8'b00110010: bin_r = 8'b00100011;  // gc: 50, bin: 35
        8'b00110110: bin_r = 8'b00100100;  // gc: 54, bin: 36
        8'b00110111: bin_r = 8'b00100101;  // gc: 55, bin: 37
        8'b00110101: bin_r = 8'b00100110;  // gc: 53, bin: 38
        8'b00110100: bin_r = 8'b00100111;  // gc: 52, bin: 39
        8'b00111100: bin_r = 8'b00101000;  // gc: 60, bin: 40
        8'b00111101: bin_r = 8'b00101001;  // gc: 61, bin: 41
        8'b00111111: bin_r = 8'b00101010;  // gc: 63, bin: 42
        8'b00111110: bin_r = 8'b00101011;  // gc: 62, bin: 43
        8'b00111010: bin_r = 8'b00101100;  // gc: 58, bin: 44
        8'b00111011: bin_r = 8'b00101101;  // gc: 59, bin: 45
        8'b00111001: bin_r = 8'b00101110;  // gc: 57, bin: 46
        8'b00111000: bin_r = 8'b00101111;  // gc: 56, bin: 47
        8'b00101000: bin_r = 8'b00110000;  // gc: 40, bin: 48
        8'b00101001: bin_r = 8'b00110001;  // gc: 41, bin: 49
        8'b00101011: bin_r = 8'b00110010;  // gc: 43, bin: 50
        8'b00101010: bin_r = 8'b00110011;  // gc: 42, bin: 51
        8'b00101110: bin_r = 8'b00110100;  // gc: 46, bin: 52
        8'b00101111: bin_r = 8'b00110101;  // gc: 47, bin: 53
        8'b00101101: bin_r = 8'b00110110;  // gc: 45, bin: 54
        8'b00101100: bin_r = 8'b00110111;  // gc: 44, bin: 55
        8'b00100100: bin_r = 8'b00111000;  // gc: 36, bin: 56
        8'b00100101: bin_r = 8'b00111001;  // gc: 37, bin: 57
        8'b00100111: bin_r = 8'b00111010;  // gc: 39, bin: 58
        8'b00100110: bin_r = 8'b00111011;  // gc: 38, bin: 59
        8'b00100010: bin_r = 8'b00111100;  // gc: 34, bin: 60
        8'b00100011: bin_r = 8'b00111101;  // gc: 35, bin: 61
        8'b00100001: bin_r = 8'b00111110;  // gc: 33, bin: 62
        8'b00100000: bin_r = 8'b00111111;  // gc: 32, bin: 63
        8'b01100000: bin_r = 8'b01000000;  // gc: 96, bin: 64
        8'b01100001: bin_r = 8'b01000001;  // gc: 97, bin: 65
        8'b01100011: bin_r = 8'b01000010;  // gc: 99, bin: 66
        8'b01100010: bin_r = 8'b01000011;  // gc: 98, bin: 67
        8'b01100110: bin_r = 8'b01000100;  // gc: 102, bin: 68
        8'b01100111: bin_r = 8'b01000101;  // gc: 103, bin: 69
        8'b01100101: bin_r = 8'b01000110;  // gc: 101, bin: 70
        8'b01100100: bin_r = 8'b01000111;  // gc: 100, bin: 71
        8'b01101100: bin_r = 8'b01001000;  // gc: 108, bin: 72
        8'b01101101: bin_r = 8'b01001001;  // gc: 109, bin: 73
        8'b01101111: bin_r = 8'b01001010;  // gc: 111, bin: 74
        8'b01101110: bin_r = 8'b01001011;  // gc: 110, bin: 75
        8'b01101010: bin_r = 8'b01001100;  // gc: 106, bin: 76
        8'b01101011: bin_r = 8'b01001101;  // gc: 107, bin: 77
        8'b01101001: bin_r = 8'b01001110;  // gc: 105, bin: 78
        8'b01101000: bin_r = 8'b01001111;  // gc: 104, bin: 79
        8'b01111000: bin_r = 8'b01010000;  // gc: 120, bin: 80
        8'b01111001: bin_r = 8'b01010001;  // gc: 121, bin: 81
        8'b01111011: bin_r = 8'b01010010;  // gc: 123, bin: 82
        8'b01111010: bin_r = 8'b01010011;  // gc: 122, bin: 83
        8'b01111110: bin_r = 8'b01010100;  // gc: 126, bin: 84
        8'b01111111: bin_r = 8'b01010101;  // gc: 127, bin: 85
        8'b01111101: bin_r = 8'b01010110;  // gc: 125, bin: 86
        8'b01111100: bin_r = 8'b01010111;  // gc: 124, bin: 87
        8'b01110100: bin_r = 8'b01011000;  // gc: 116, bin: 88
        8'b01110101: bin_r = 8'b01011001;  // gc: 117, bin: 89
        8'b01110111: bin_r = 8'b01011010;  // gc: 119, bin: 90
        8'b01110110: bin_r = 8'b01011011;  // gc: 118, bin: 91
        8'b01110010: bin_r = 8'b01011100;  // gc: 114, bin: 92
        8'b01110011: bin_r = 8'b01011101;  // gc: 115, bin: 93
        8'b01110001: bin_r = 8'b01011110;  // gc: 113, bin: 94
        8'b01110000: bin_r = 8'b01011111;  // gc: 112, bin: 95
        8'b01010000: bin_r = 8'b01100000;  // gc: 80, bin: 96
        8'b01010001: bin_r = 8'b01100001;  // gc: 81, bin: 97
        8'b01010011: bin_r = 8'b01100010;  // gc: 83, bin: 98
        8'b01010010: bin_r = 8'b01100011;  // gc: 82, bin: 99
        8'b01010110: bin_r = 8'b01100100;  // gc: 86, bin: 100
        8'b01010111: bin_r = 8'b01100101;  // gc: 87, bin: 101
        8'b01010101: bin_r = 8'b01100110;  // gc: 85, bin: 102
        8'b01010100: bin_r = 8'b01100111;  // gc: 84, bin: 103
        8'b01011100: bin_r = 8'b01101000;  // gc: 92, bin: 104
        8'b01011101: bin_r = 8'b01101001;  // gc: 93, bin: 105
        8'b01011111: bin_r = 8'b01101010;  // gc: 95, bin: 106
        8'b01011110: bin_r = 8'b01101011;  // gc: 94, bin: 107
        8'b01011010: bin_r = 8'b01101100;  // gc: 90, bin: 108
        8'b01011011: bin_r = 8'b01101101;  // gc: 91, bin: 109
        8'b01011001: bin_r = 8'b01101110;  // gc: 89, bin: 110
        8'b01011000: bin_r = 8'b01101111;  // gc: 88, bin: 111
        8'b01001000: bin_r = 8'b01110000;  // gc: 72, bin: 112
        8'b01001001: bin_r = 8'b01110001;  // gc: 73, bin: 113
        8'b01001011: bin_r = 8'b01110010;  // gc: 75, bin: 114
        8'b01001010: bin_r = 8'b01110011;  // gc: 74, bin: 115
        8'b01001110: bin_r = 8'b01110100;  // gc: 78, bin: 116
        8'b01001111: bin_r = 8'b01110101;  // gc: 79, bin: 117
        8'b01001101: bin_r = 8'b01110110;  // gc: 77, bin: 118
        8'b01001100: bin_r = 8'b01110111;  // gc: 76, bin: 119
        8'b01000100: bin_r = 8'b01111000;  // gc: 68, bin: 120
        8'b01000101: bin_r = 8'b01111001;  // gc: 69, bin: 121
        8'b01000111: bin_r = 8'b01111010;  // gc: 71, bin: 122
        8'b01000110: bin_r = 8'b01111011;  // gc: 70, bin: 123
        8'b01000010: bin_r = 8'b01111100;  // gc: 66, bin: 124
        8'b01000011: bin_r = 8'b01111101;  // gc: 67, bin: 125
        8'b01000001: bin_r = 8'b01111110;  // gc: 65, bin: 126
        8'b01000000: bin_r = 8'b01111111;  // gc: 64, bin: 127
        8'b11000000: bin_r = 8'b10000000;  // gc: 192, bin: 128
        8'b11000001: bin_r = 8'b10000001;  // gc: 193, bin: 129
        8'b11000011: bin_r = 8'b10000010;  // gc: 195, bin: 130
        8'b11000010: bin_r = 8'b10000011;  // gc: 194, bin: 131
        8'b11000110: bin_r = 8'b10000100;  // gc: 198, bin: 132
        8'b11000111: bin_r = 8'b10000101;  // gc: 199, bin: 133
        8'b11000101: bin_r = 8'b10000110;  // gc: 197, bin: 134
        8'b11000100: bin_r = 8'b10000111;  // gc: 196, bin: 135
        8'b11001100: bin_r = 8'b10001000;  // gc: 204, bin: 136
        8'b11001101: bin_r = 8'b10001001;  // gc: 205, bin: 137
        8'b11001111: bin_r = 8'b10001010;  // gc: 207, bin: 138
        8'b11001110: bin_r = 8'b10001011;  // gc: 206, bin: 139
        8'b11001010: bin_r = 8'b10001100;  // gc: 202, bin: 140
        8'b11001011: bin_r = 8'b10001101;  // gc: 203, bin: 141
        8'b11001001: bin_r = 8'b10001110;  // gc: 201, bin: 142
        8'b11001000: bin_r = 8'b10001111;  // gc: 200, bin: 143
        8'b11011000: bin_r = 8'b10010000;  // gc: 216, bin: 144
        8'b11011001: bin_r = 8'b10010001;  // gc: 217, bin: 145
        8'b11011011: bin_r = 8'b10010010;  // gc: 219, bin: 146
        8'b11011010: bin_r = 8'b10010011;  // gc: 218, bin: 147
        8'b11011110: bin_r = 8'b10010100;  // gc: 222, bin: 148
        8'b11011111: bin_r = 8'b10010101;  // gc: 223, bin: 149
        8'b11011101: bin_r = 8'b10010110;  // gc: 221, bin: 150
        8'b11011100: bin_r = 8'b10010111;  // gc: 220, bin: 151
        8'b11010100: bin_r = 8'b10011000;  // gc: 212, bin: 152
        8'b11010101: bin_r = 8'b10011001;  // gc: 213, bin: 153
        8'b11010111: bin_r = 8'b10011010;  // gc: 215, bin: 154
        8'b11010110: bin_r = 8'b10011011;  // gc: 214, bin: 155
        8'b11010010: bin_r = 8'b10011100;  // gc: 210, bin: 156
        8'b11010011: bin_r = 8'b10011101;  // gc: 211, bin: 157
        8'b11010001: bin_r = 8'b10011110;  // gc: 209, bin: 158
        8'b11010000: bin_r = 8'b10011111;  // gc: 208, bin: 159
        8'b11110000: bin_r = 8'b10100000;  // gc: 240, bin: 160
        8'b11110001: bin_r = 8'b10100001;  // gc: 241, bin: 161
        8'b11110011: bin_r = 8'b10100010;  // gc: 243, bin: 162
        8'b11110010: bin_r = 8'b10100011;  // gc: 242, bin: 163
        8'b11110110: bin_r = 8'b10100100;  // gc: 246, bin: 164
        8'b11110111: bin_r = 8'b10100101;  // gc: 247, bin: 165
        8'b11110101: bin_r = 8'b10100110;  // gc: 245, bin: 166
        8'b11110100: bin_r = 8'b10100111;  // gc: 244, bin: 167
        8'b11111100: bin_r = 8'b10101000;  // gc: 252, bin: 168
        8'b11111101: bin_r = 8'b10101001;  // gc: 253, bin: 169
        8'b11111111: bin_r = 8'b10101010;  // gc: 255, bin: 170
        8'b11111110: bin_r = 8'b10101011;  // gc: 254, bin: 171
        8'b11111010: bin_r = 8'b10101100;  // gc: 250, bin: 172
        8'b11111011: bin_r = 8'b10101101;  // gc: 251, bin: 173
        8'b11111001: bin_r = 8'b10101110;  // gc: 249, bin: 174
        8'b11111000: bin_r = 8'b10101111;  // gc: 248, bin: 175
        8'b11101000: bin_r = 8'b10110000;  // gc: 232, bin: 176
        8'b11101001: bin_r = 8'b10110001;  // gc: 233, bin: 177
        8'b11101011: bin_r = 8'b10110010;  // gc: 235, bin: 178
        8'b11101010: bin_r = 8'b10110011;  // gc: 234, bin: 179
        8'b11101110: bin_r = 8'b10110100;  // gc: 238, bin: 180
        8'b11101111: bin_r = 8'b10110101;  // gc: 239, bin: 181
        8'b11101101: bin_r = 8'b10110110;  // gc: 237, bin: 182
        8'b11101100: bin_r = 8'b10110111;  // gc: 236, bin: 183
        8'b11100100: bin_r = 8'b10111000;  // gc: 228, bin: 184
        8'b11100101: bin_r = 8'b10111001;  // gc: 229, bin: 185
        8'b11100111: bin_r = 8'b10111010;  // gc: 231, bin: 186
        8'b11100110: bin_r = 8'b10111011;  // gc: 230, bin: 187
        8'b11100010: bin_r = 8'b10111100;  // gc: 226, bin: 188
        8'b11100011: bin_r = 8'b10111101;  // gc: 227, bin: 189
        8'b11100001: bin_r = 8'b10111110;  // gc: 225, bin: 190
        8'b11100000: bin_r = 8'b10111111;  // gc: 224, bin: 191
        8'b10100000: bin_r = 8'b11000000;  // gc: 160, bin: 192
        8'b10100001: bin_r = 8'b11000001;  // gc: 161, bin: 193
        8'b10100011: bin_r = 8'b11000010;  // gc: 163, bin: 194
        8'b10100010: bin_r = 8'b11000011;  // gc: 162, bin: 195
        8'b10100110: bin_r = 8'b11000100;  // gc: 166, bin: 196
        8'b10100111: bin_r = 8'b11000101;  // gc: 167, bin: 197
        8'b10100101: bin_r = 8'b11000110;  // gc: 165, bin: 198
        8'b10100100: bin_r = 8'b11000111;  // gc: 164, bin: 199
        8'b10101100: bin_r = 8'b11001000;  // gc: 172, bin: 200
        8'b10101101: bin_r = 8'b11001001;  // gc: 173, bin: 201
        8'b10101111: bin_r = 8'b11001010;  // gc: 175, bin: 202
        8'b10101110: bin_r = 8'b11001011;  // gc: 174, bin: 203
        8'b10101010: bin_r = 8'b11001100;  // gc: 170, bin: 204
        8'b10101011: bin_r = 8'b11001101;  // gc: 171, bin: 205
        8'b10101001: bin_r = 8'b11001110;  // gc: 169, bin: 206
        8'b10101000: bin_r = 8'b11001111;  // gc: 168, bin: 207
        8'b10111000: bin_r = 8'b11010000;  // gc: 184, bin: 208
        8'b10111001: bin_r = 8'b11010001;  // gc: 185, bin: 209
        8'b10111011: bin_r = 8'b11010010;  // gc: 187, bin: 210
        8'b10111010: bin_r = 8'b11010011;  // gc: 186, bin: 211
        8'b10111110: bin_r = 8'b11010100;  // gc: 190, bin: 212
        8'b10111111: bin_r = 8'b11010101;  // gc: 191, bin: 213
        8'b10111101: bin_r = 8'b11010110;  // gc: 189, bin: 214
        8'b10111100: bin_r = 8'b11010111;  // gc: 188, bin: 215
        8'b10110100: bin_r = 8'b11011000;  // gc: 180, bin: 216
        8'b10110101: bin_r = 8'b11011001;  // gc: 181, bin: 217
        8'b10110111: bin_r = 8'b11011010;  // gc: 183, bin: 218
        8'b10110110: bin_r = 8'b11011011;  // gc: 182, bin: 219
        8'b10110010: bin_r = 8'b11011100;  // gc: 178, bin: 220
        8'b10110011: bin_r = 8'b11011101;  // gc: 179, bin: 221
        8'b10110001: bin_r = 8'b11011110;  // gc: 177, bin: 222
        8'b10110000: bin_r = 8'b11011111;  // gc: 176, bin: 223
        8'b10010000: bin_r = 8'b11100000;  // gc: 144, bin: 224
        8'b10010001: bin_r = 8'b11100001;  // gc: 145, bin: 225
        8'b10010011: bin_r = 8'b11100010;  // gc: 147, bin: 226
        8'b10010010: bin_r = 8'b11100011;  // gc: 146, bin: 227
        8'b10010110: bin_r = 8'b11100100;  // gc: 150, bin: 228
        8'b10010111: bin_r = 8'b11100101;  // gc: 151, bin: 229
        8'b10010101: bin_r = 8'b11100110;  // gc: 149, bin: 230
        8'b10010100: bin_r = 8'b11100111;  // gc: 148, bin: 231
        8'b10011100: bin_r = 8'b11101000;  // gc: 156, bin: 232
        8'b10011101: bin_r = 8'b11101001;  // gc: 157, bin: 233
        8'b10011111: bin_r = 8'b11101010;  // gc: 159, bin: 234
        8'b10011110: bin_r = 8'b11101011;  // gc: 158, bin: 235
        8'b10011010: bin_r = 8'b11101100;  // gc: 154, bin: 236
        8'b10011011: bin_r = 8'b11101101;  // gc: 155, bin: 237
        8'b10011001: bin_r = 8'b11101110;  // gc: 153, bin: 238
        8'b10011000: bin_r = 8'b11101111;  // gc: 152, bin: 239
        8'b10001000: bin_r = 8'b11110000;  // gc: 136, bin: 240
        8'b10001001: bin_r = 8'b11110001;  // gc: 137, bin: 241
        8'b10001011: bin_r = 8'b11110010;  // gc: 139, bin: 242
        8'b10001010: bin_r = 8'b11110011;  // gc: 138, bin: 243
        8'b10001110: bin_r = 8'b11110100;  // gc: 142, bin: 244
        8'b10001111: bin_r = 8'b11110101;  // gc: 143, bin: 245
        8'b10001101: bin_r = 8'b11110110;  // gc: 141, bin: 246
        8'b10001100: bin_r = 8'b11110111;  // gc: 140, bin: 247
        8'b10000100: bin_r = 8'b11111000;  // gc: 132, bin: 248
        8'b10000101: bin_r = 8'b11111001;  // gc: 133, bin: 249
        8'b10000111: bin_r = 8'b11111010;  // gc: 135, bin: 250
        8'b10000110: bin_r = 8'b11111011;  // gc: 134, bin: 251
        8'b10000010: bin_r = 8'b11111100;  // gc: 130, bin: 252
        8'b10000011: bin_r = 8'b11111101;  // gc: 131, bin: 253
        8'b10000001: bin_r = 8'b11111110;  // gc: 129, bin: 254
        8'b10000000: bin_r = 8'b11111111;  // gc: 128, bin: 255
        default: bin_r = 8'd0; // Fully described
    endcase
end

endmodule

